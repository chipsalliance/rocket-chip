`ifndef CONST_VH
`define CONST_VH

`define MEM_ADDR_BITS 34
`define MEM_DATA_BITS 128
`define MEM_TAG_BITS 10

`endif // CONST_VH
